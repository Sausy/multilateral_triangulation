// test_programm.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module test_programm (
		input  wire       clk_clk,                    //       clk.clk
		input  wire       reset_reset_n,              //     reset.reset_n
		input  wire       spislave0_ispi_in,          // spislave0.ispi_in
		input  wire [7:0] spislave0_ispi_send_byte,   //          .ispi_send_byte
		input  wire       spislave0_ispi_ss_n,        //          .ispi_ss_n
		output wire       spislave0_ospi_inc_wraddr,  //          .ospi_inc_wraddr
		output wire       spislave0_ospi_out,         //          .ospi_out
		output wire [4:0] spislave0_ospi_periph_slct, //          .ospi_periph_slct
		output wire [7:0] spislave0_ospi_rcv_byte,    //          .ospi_rcv_byte
		output wire [7:0] spislave0_ospi_rcv_cmd,     //          .ospi_rcv_cmd
		output wire       spislave0_ospi_write_sig    //          .ospi_write_sig
	);

	SPISlave spislave_0 (
		.clk              (clk_clk),                    //       clock.clk
		.iSPI_IN          (spislave0_ispi_in),          // conduit_end.ispi_in
		.iSPI_SEND_BYTE   (spislave0_ispi_send_byte),   //            .ispi_send_byte
		.iSPI_SS_n        (spislave0_ispi_ss_n),        //            .ispi_ss_n
		.oSPI_INC_WRADDR  (spislave0_ospi_inc_wraddr),  //            .ospi_inc_wraddr
		.oSPI_OUT         (spislave0_ospi_out),         //            .ospi_out
		.oSPI_PERIPH_SLCT (spislave0_ospi_periph_slct), //            .ospi_periph_slct
		.oSPI_RCV_BYTE    (spislave0_ospi_rcv_byte),    //            .ospi_rcv_byte
		.oSPI_RCV_CMD     (spislave0_ospi_rcv_cmd),     //            .ospi_rcv_cmd
		.oSPI_WRITE_SIG   (spislave0_ospi_write_sig)    //            .ospi_write_sig
	);

endmodule
