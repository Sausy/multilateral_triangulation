// soc_system.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                                       //                           clk.clk
		output wire        clock_divider_0_conduit_end_out_clk,           //   clock_divider_0_conduit_end.out_clk
		input  wire [1:0]  fpga_key_input_export,                         //                fpga_key_input.export
		output wire [7:0]  fpga_led_output_export,                        //               fpga_led_output.export
		output wire [14:0] hps_ddr_mem_a,                                 //                       hps_ddr.mem_a
		output wire [2:0]  hps_ddr_mem_ba,                                //                              .mem_ba
		output wire        hps_ddr_mem_ck,                                //                              .mem_ck
		output wire        hps_ddr_mem_ck_n,                              //                              .mem_ck_n
		output wire        hps_ddr_mem_cke,                               //                              .mem_cke
		output wire        hps_ddr_mem_cs_n,                              //                              .mem_cs_n
		output wire        hps_ddr_mem_ras_n,                             //                              .mem_ras_n
		output wire        hps_ddr_mem_cas_n,                             //                              .mem_cas_n
		output wire        hps_ddr_mem_we_n,                              //                              .mem_we_n
		output wire        hps_ddr_mem_reset_n,                           //                              .mem_reset_n
		inout  wire [31:0] hps_ddr_mem_dq,                                //                              .mem_dq
		inout  wire [3:0]  hps_ddr_mem_dqs,                               //                              .mem_dqs
		inout  wire [3:0]  hps_ddr_mem_dqs_n,                             //                              .mem_dqs_n
		output wire        hps_ddr_mem_odt,                               //                              .mem_odt
		output wire [3:0]  hps_ddr_mem_dm,                                //                              .mem_dm
		input  wire        hps_ddr_oct_rzqin,                             //                              .oct_rzqin
		output wire [66:0] hps_h2f_loan_io_in,                            //               hps_h2f_loan_io.in
		input  wire [66:0] hps_h2f_loan_io_out,                           //                              .out
		input  wire [66:0] hps_h2f_loan_io_oe,                            //                              .oe
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,               //                        hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,                 //                              .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,                 //                              .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,                 //                              .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,                 //                              .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,                 //                              .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,                 //                              .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,                  //                              .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,               //                              .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,               //                              .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,               //                              .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,                 //                              .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,                 //                              .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,                 //                              .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                   //                              .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                    //                              .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                    //                              .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,                   //                              .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                    //                              .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                    //                              .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                    //                              .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                    //                              .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                    //                              .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                    //                              .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                    //                              .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                    //                              .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                    //                              .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                    //                              .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                   //                              .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                   //                              .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                   //                              .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                   //                              .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,                   //                              .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                   //                              .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,                   //                              .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,                   //                              .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,                //                              .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,                //                              .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,                //                              .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,                //                              .hps_io_gpio_inst_GPIO61
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO40,              //                              .hps_io_gpio_inst_LOANIO40
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO51,              //                              .hps_io_gpio_inst_LOANIO51
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO52,              //                              .hps_io_gpio_inst_LOANIO52
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO54,              //                              .hps_io_gpio_inst_LOANIO54
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO64,              //                              .hps_io_gpio_inst_LOANIO64
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO65,              //                              .hps_io_gpio_inst_LOANIO65
		input  wire [3:0]  id_switch0_sw,                                 //                    id_switch0.sw
		output wire        piezo_controller_piezo_enable_export,          // piezo_controller_piezo_enable.export
		input  wire        piezo_controller_piezo_enable_piezo_enable_in, //                              .piezo_enable_in
		output wire [60:0] piezo_controller_piezo_out_export,             //    piezo_controller_piezo_out.export
		output wire [2:0]  piezo_controller_piezo_status_export,          // piezo_controller_piezo_status.export
		input  wire        ptp_piezo_interface0_piezo_interface_in,       //          ptp_piezo_interface0.piezo_interface_in
		output wire        ptp_piezo_interface0_piezo_interface_out,      //                              .piezo_interface_out
		input  wire        reset_reset_n,                                 //                         reset.reset_n
		input  wire        rtc_0_conduit_end_event_trigger,               //             rtc_0_conduit_end.event_trigger
		output wire        rtc_0_conduit_end_piezo_enable,                //                              .piezo_enable
		input  wire        rtc_0_conduit_end_event_trigger2               //                              .event_trigger2
	);

	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                      // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                        // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                        // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                       // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                       // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                        // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                          // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                      // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                       // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                       // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                       // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                       // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                        // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                      // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                      // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                         // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                       // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                       // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                       // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                      // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                       // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                       // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                        // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                         // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                       // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                       // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                      // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                       // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_realtime_clock_controll_0_avalon_slave_readdata;    // realtime_clock_controll_0:avalon_slave_readdata -> mm_interconnect_0:realtime_clock_controll_0_avalon_slave_readdata
	wire         mm_interconnect_0_realtime_clock_controll_0_avalon_slave_waitrequest; // realtime_clock_controll_0:avalon_slave_waitrequest -> mm_interconnect_0:realtime_clock_controll_0_avalon_slave_waitrequest
	wire  [15:0] mm_interconnect_0_realtime_clock_controll_0_avalon_slave_address;     // mm_interconnect_0:realtime_clock_controll_0_avalon_slave_address -> realtime_clock_controll_0:avalon_slave_address
	wire         mm_interconnect_0_realtime_clock_controll_0_avalon_slave_read;        // mm_interconnect_0:realtime_clock_controll_0_avalon_slave_read -> realtime_clock_controll_0:avalon_slave_read
	wire         mm_interconnect_0_realtime_clock_controll_0_avalon_slave_write;       // mm_interconnect_0:realtime_clock_controll_0_avalon_slave_write -> realtime_clock_controll_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_realtime_clock_controll_0_avalon_slave_writedata;   // mm_interconnect_0:realtime_clock_controll_0_avalon_slave_writedata -> realtime_clock_controll_0:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_ptp_simple_us_0_avalon_slave_readdata;              // ptp_simple_us_0:avalon_slave_readdata -> mm_interconnect_0:ptp_simple_us_0_avalon_slave_readdata
	wire         mm_interconnect_0_ptp_simple_us_0_avalon_slave_waitrequest;           // ptp_simple_us_0:avalon_slave_waitrequest -> mm_interconnect_0:ptp_simple_us_0_avalon_slave_waitrequest
	wire  [15:0] mm_interconnect_0_ptp_simple_us_0_avalon_slave_address;               // mm_interconnect_0:ptp_simple_us_0_avalon_slave_address -> ptp_simple_us_0:avalon_slave_address
	wire         mm_interconnect_0_ptp_simple_us_0_avalon_slave_read;                  // mm_interconnect_0:ptp_simple_us_0_avalon_slave_read -> ptp_simple_us_0:avalon_slave_read
	wire         mm_interconnect_0_ptp_simple_us_0_avalon_slave_write;                 // mm_interconnect_0:ptp_simple_us_0_avalon_slave_write -> ptp_simple_us_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_ptp_simple_us_0_avalon_slave_writedata;             // mm_interconnect_0:ptp_simple_us_0_avalon_slave_writedata -> ptp_simple_us_0:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_id_switch_0_avalon_slave_readdata;                  // id_switch_0:avalon_slave_readdata -> mm_interconnect_0:id_switch_0_avalon_slave_readdata
	wire         mm_interconnect_0_id_switch_0_avalon_slave_waitrequest;               // id_switch_0:avalon_slave_waitrequest -> mm_interconnect_0:id_switch_0_avalon_slave_waitrequest
	wire  [15:0] mm_interconnect_0_id_switch_0_avalon_slave_address;                   // mm_interconnect_0:id_switch_0_avalon_slave_address -> id_switch_0:avalon_slave_address
	wire         mm_interconnect_0_id_switch_0_avalon_slave_read;                      // mm_interconnect_0:id_switch_0_avalon_slave_read -> id_switch_0:avalon_slave_read
	wire         mm_interconnect_0_id_switch_0_avalon_slave_write;                     // mm_interconnect_0:id_switch_0_avalon_slave_write -> id_switch_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_id_switch_0_avalon_slave_writedata;                 // mm_interconnect_0:id_switch_0_avalon_slave_writedata -> id_switch_0:avalon_slave_writedata
	wire         mm_interconnect_0_fpga_key_s1_chipselect;                             // mm_interconnect_0:fpga_key_s1_chipselect -> fpga_key:chipselect
	wire  [31:0] mm_interconnect_0_fpga_key_s1_readdata;                               // fpga_key:readdata -> mm_interconnect_0:fpga_key_s1_readdata
	wire   [1:0] mm_interconnect_0_fpga_key_s1_address;                                // mm_interconnect_0:fpga_key_s1_address -> fpga_key:address
	wire         mm_interconnect_0_fpga_key_s1_write;                                  // mm_interconnect_0:fpga_key_s1_write -> fpga_key:write_n
	wire  [31:0] mm_interconnect_0_fpga_key_s1_writedata;                              // mm_interconnect_0:fpga_key_s1_writedata -> fpga_key:writedata
	wire         mm_interconnect_0_fpga_led_s1_chipselect;                             // mm_interconnect_0:fpga_led_s1_chipselect -> fpga_led:chipselect
	wire  [31:0] mm_interconnect_0_fpga_led_s1_readdata;                               // fpga_led:readdata -> mm_interconnect_0:fpga_led_s1_readdata
	wire   [2:0] mm_interconnect_0_fpga_led_s1_address;                                // mm_interconnect_0:fpga_led_s1_address -> fpga_led:address
	wire         mm_interconnect_0_fpga_led_s1_write;                                  // mm_interconnect_0:fpga_led_s1_write -> fpga_led:write_n
	wire  [31:0] mm_interconnect_0_fpga_led_s1_writedata;                              // mm_interconnect_0:fpga_led_s1_writedata -> fpga_led:writedata
	wire  [15:0] mm_interconnect_0_piezo_controller_0_s1_readdata;                     // piezo_controller_0:AVS_ReadData -> mm_interconnect_0:piezo_controller_0_s1_readdata
	wire   [7:0] mm_interconnect_0_piezo_controller_0_s1_address;                      // mm_interconnect_0:piezo_controller_0_s1_address -> piezo_controller_0:AVS_Address
	wire         mm_interconnect_0_piezo_controller_0_s1_read;                         // mm_interconnect_0:piezo_controller_0_s1_read -> piezo_controller_0:AVS_Read
	wire         mm_interconnect_0_piezo_controller_0_s1_write;                        // mm_interconnect_0:piezo_controller_0_s1_write -> piezo_controller_0:AVS_Write
	wire  [15:0] mm_interconnect_0_piezo_controller_0_s1_writedata;                    // mm_interconnect_0:piezo_controller_0_s1_writedata -> piezo_controller_0:AVS_WriteData
	wire         irq_mapper_receiver0_irq;                                             // fpga_key:irq -> irq_mapper:receiver0_irq
	wire  [31:0] hps_0_f2h_irq0_irq;                                                   // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                                   // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [clock_divider_0:reset, id_switch_0:reset, mm_interconnect_0:realtime_clock_controll_0_reset_reset_bridge_in_reset_reset, ptp_simple_us_0:reset, realtime_clock_controll_0:reset]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [fpga_key:reset_n, fpga_led:reset_n, mm_interconnect_0:fpga_key_reset_reset_bridge_in_reset_reset, piezo_controller_0:reset_n]
	wire         hps_0_h2f_reset_reset;                                                // hps_0:h2f_rst_n -> [rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire         rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	clock_divider clock_divider_0 (
		.clock   (clk_clk),                             //  clock_sink.clk
		.reset   (rst_controller_reset_out_reset),      //       reset.reset
		.out_clk (clock_divider_0_conduit_end_out_clk)  // conduit_end.out_clk
	);

	soc_system_fpga_key fpga_key (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_fpga_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fpga_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fpga_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fpga_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fpga_key_s1_readdata),   //                    .readdata
		.in_port    (fpga_key_input_export),                    // external_connection.export
		.irq        (irq_mapper_receiver0_irq)                  //                 irq.irq
	);

	soc_system_fpga_led fpga_led (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_fpga_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fpga_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fpga_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fpga_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fpga_led_s1_readdata),   //                    .readdata
		.out_port   (fpga_led_output_export)                    // external_connection.export
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_loan_in               (hps_h2f_loan_io_in),               //       h2f_loan_io.in
		.h2f_loan_out              (hps_h2f_loan_io_out),              //                  .out
		.h2f_loan_oe               (hps_h2f_loan_io_oe),               //                  .oe
		.mem_a                     (hps_ddr_mem_a),                    //            memory.mem_a
		.mem_ba                    (hps_ddr_mem_ba),                   //                  .mem_ba
		.mem_ck                    (hps_ddr_mem_ck),                   //                  .mem_ck
		.mem_ck_n                  (hps_ddr_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                   (hps_ddr_mem_cke),                  //                  .mem_cke
		.mem_cs_n                  (hps_ddr_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                 (hps_ddr_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                 (hps_ddr_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                  (hps_ddr_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n               (hps_ddr_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                    (hps_ddr_mem_dq),                   //                  .mem_dq
		.mem_dqs                   (hps_ddr_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                 (hps_ddr_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                   (hps_ddr_mem_odt),                  //                  .mem_odt
		.mem_dm                    (hps_ddr_mem_dm),                   //                  .mem_dm
		.oct_rzqin                 (hps_ddr_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK  (hps_io_hps_io_emac1_inst_TX_CLK),  //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0    (hps_io_hps_io_emac1_inst_TXD0),    //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1    (hps_io_hps_io_emac1_inst_TXD1),    //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2    (hps_io_hps_io_emac1_inst_TXD2),    //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3    (hps_io_hps_io_emac1_inst_TXD3),    //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0    (hps_io_hps_io_emac1_inst_RXD0),    //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO    (hps_io_hps_io_emac1_inst_MDIO),    //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC     (hps_io_hps_io_emac1_inst_MDC),     //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL  (hps_io_hps_io_emac1_inst_RX_CTL),  //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL  (hps_io_hps_io_emac1_inst_TX_CTL),  //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK  (hps_io_hps_io_emac1_inst_RX_CLK),  //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1    (hps_io_hps_io_emac1_inst_RXD1),    //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2    (hps_io_hps_io_emac1_inst_RXD2),    //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3    (hps_io_hps_io_emac1_inst_RXD3),    //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD      (hps_io_hps_io_sdio_inst_CMD),      //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_io_hps_io_sdio_inst_D0),       //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_io_hps_io_sdio_inst_D1),       //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_io_hps_io_sdio_inst_CLK),      //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_io_hps_io_sdio_inst_D2),       //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_io_hps_io_sdio_inst_D3),       //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0       (hps_io_hps_io_usb1_inst_D0),       //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1       (hps_io_hps_io_usb1_inst_D1),       //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2       (hps_io_hps_io_usb1_inst_D2),       //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3       (hps_io_hps_io_usb1_inst_D3),       //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4       (hps_io_hps_io_usb1_inst_D4),       //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5       (hps_io_hps_io_usb1_inst_D5),       //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6       (hps_io_hps_io_usb1_inst_D6),       //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7       (hps_io_hps_io_usb1_inst_D7),       //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK      (hps_io_hps_io_usb1_inst_CLK),      //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP      (hps_io_hps_io_usb1_inst_STP),      //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR      (hps_io_hps_io_usb1_inst_DIR),      //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT      (hps_io_hps_io_usb1_inst_NXT),      //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX      (hps_io_hps_io_uart0_inst_RX),      //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX      (hps_io_hps_io_uart0_inst_TX),      //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA      (hps_io_hps_io_i2c0_inst_SDA),      //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL      (hps_io_hps_io_i2c0_inst_SCL),      //                  .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO09   (hps_io_hps_io_gpio_inst_GPIO09),   //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35   (hps_io_hps_io_gpio_inst_GPIO35),   //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO53   (hps_io_hps_io_gpio_inst_GPIO53),   //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO61   (hps_io_hps_io_gpio_inst_GPIO61),   //                  .hps_io_gpio_inst_GPIO61
		.hps_io_gpio_inst_LOANIO40 (hps_io_hps_io_gpio_inst_LOANIO40), //                  .hps_io_gpio_inst_LOANIO40
		.hps_io_gpio_inst_LOANIO51 (hps_io_hps_io_gpio_inst_LOANIO51), //                  .hps_io_gpio_inst_LOANIO51
		.hps_io_gpio_inst_LOANIO52 (hps_io_hps_io_gpio_inst_LOANIO52), //                  .hps_io_gpio_inst_LOANIO52
		.hps_io_gpio_inst_LOANIO54 (hps_io_hps_io_gpio_inst_LOANIO54), //                  .hps_io_gpio_inst_LOANIO54
		.hps_io_gpio_inst_LOANIO64 (hps_io_hps_io_gpio_inst_LOANIO64), //                  .hps_io_gpio_inst_LOANIO64
		.hps_io_gpio_inst_LOANIO65 (hps_io_hps_io_gpio_inst_LOANIO65), //                  .hps_io_gpio_inst_LOANIO65
		.h2f_rst_n                 (hps_0_h2f_reset_reset),            //         h2f_reset.reset_n
		.h2f_lw_axi_clk            (clk_clk),                          //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID               (hps_0_h2f_lw_axi_master_awid),     // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR             (hps_0_h2f_lw_axi_master_awaddr),   //                  .awaddr
		.h2f_lw_AWLEN              (hps_0_h2f_lw_axi_master_awlen),    //                  .awlen
		.h2f_lw_AWSIZE             (hps_0_h2f_lw_axi_master_awsize),   //                  .awsize
		.h2f_lw_AWBURST            (hps_0_h2f_lw_axi_master_awburst),  //                  .awburst
		.h2f_lw_AWLOCK             (hps_0_h2f_lw_axi_master_awlock),   //                  .awlock
		.h2f_lw_AWCACHE            (hps_0_h2f_lw_axi_master_awcache),  //                  .awcache
		.h2f_lw_AWPROT             (hps_0_h2f_lw_axi_master_awprot),   //                  .awprot
		.h2f_lw_AWVALID            (hps_0_h2f_lw_axi_master_awvalid),  //                  .awvalid
		.h2f_lw_AWREADY            (hps_0_h2f_lw_axi_master_awready),  //                  .awready
		.h2f_lw_WID                (hps_0_h2f_lw_axi_master_wid),      //                  .wid
		.h2f_lw_WDATA              (hps_0_h2f_lw_axi_master_wdata),    //                  .wdata
		.h2f_lw_WSTRB              (hps_0_h2f_lw_axi_master_wstrb),    //                  .wstrb
		.h2f_lw_WLAST              (hps_0_h2f_lw_axi_master_wlast),    //                  .wlast
		.h2f_lw_WVALID             (hps_0_h2f_lw_axi_master_wvalid),   //                  .wvalid
		.h2f_lw_WREADY             (hps_0_h2f_lw_axi_master_wready),   //                  .wready
		.h2f_lw_BID                (hps_0_h2f_lw_axi_master_bid),      //                  .bid
		.h2f_lw_BRESP              (hps_0_h2f_lw_axi_master_bresp),    //                  .bresp
		.h2f_lw_BVALID             (hps_0_h2f_lw_axi_master_bvalid),   //                  .bvalid
		.h2f_lw_BREADY             (hps_0_h2f_lw_axi_master_bready),   //                  .bready
		.h2f_lw_ARID               (hps_0_h2f_lw_axi_master_arid),     //                  .arid
		.h2f_lw_ARADDR             (hps_0_h2f_lw_axi_master_araddr),   //                  .araddr
		.h2f_lw_ARLEN              (hps_0_h2f_lw_axi_master_arlen),    //                  .arlen
		.h2f_lw_ARSIZE             (hps_0_h2f_lw_axi_master_arsize),   //                  .arsize
		.h2f_lw_ARBURST            (hps_0_h2f_lw_axi_master_arburst),  //                  .arburst
		.h2f_lw_ARLOCK             (hps_0_h2f_lw_axi_master_arlock),   //                  .arlock
		.h2f_lw_ARCACHE            (hps_0_h2f_lw_axi_master_arcache),  //                  .arcache
		.h2f_lw_ARPROT             (hps_0_h2f_lw_axi_master_arprot),   //                  .arprot
		.h2f_lw_ARVALID            (hps_0_h2f_lw_axi_master_arvalid),  //                  .arvalid
		.h2f_lw_ARREADY            (hps_0_h2f_lw_axi_master_arready),  //                  .arready
		.h2f_lw_RID                (hps_0_h2f_lw_axi_master_rid),      //                  .rid
		.h2f_lw_RDATA              (hps_0_h2f_lw_axi_master_rdata),    //                  .rdata
		.h2f_lw_RRESP              (hps_0_h2f_lw_axi_master_rresp),    //                  .rresp
		.h2f_lw_RLAST              (hps_0_h2f_lw_axi_master_rlast),    //                  .rlast
		.h2f_lw_RVALID             (hps_0_h2f_lw_axi_master_rvalid),   //                  .rvalid
		.h2f_lw_RREADY             (hps_0_h2f_lw_axi_master_rready),   //                  .rready
		.f2h_irq_p0                (hps_0_f2h_irq0_irq),               //          f2h_irq0.irq
		.f2h_irq_p1                (hps_0_f2h_irq1_irq)                //          f2h_irq1.irq
	);

	id_switch id_switch_0 (
		.reset                    (rst_controller_reset_out_reset),                         //        reset.reset
		.avalon_slave_address     (mm_interconnect_0_id_switch_0_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_write       (mm_interconnect_0_id_switch_0_avalon_slave_write),       //             .write
		.avalon_slave_writedata   (mm_interconnect_0_id_switch_0_avalon_slave_writedata),   //             .writedata
		.avalon_slave_read        (mm_interconnect_0_id_switch_0_avalon_slave_read),        //             .read
		.avalon_slave_readdata    (mm_interconnect_0_id_switch_0_avalon_slave_readdata),    //             .readdata
		.avalon_slave_waitrequest (mm_interconnect_0_id_switch_0_avalon_slave_waitrequest), //             .waitrequest
		.sw                       (id_switch0_sw),                                          //  conduit_end.sw
		.clock                    (clk_clk)                                                 //        clock.clk
	);

	piezo_controller #(
		.piezo_count (61)
	) piezo_controller_0 (
		.clk             (clk_clk),                                           //          clk.clk
		.reset_n         (~rst_controller_001_reset_out_reset),               //        reset.reset_n
		.AVS_Address     (mm_interconnect_0_piezo_controller_0_s1_address),   //           s1.address
		.AVS_Read        (mm_interconnect_0_piezo_controller_0_s1_read),      //             .read
		.AVS_ReadData    (mm_interconnect_0_piezo_controller_0_s1_readdata),  //             .readdata
		.AVS_Write       (mm_interconnect_0_piezo_controller_0_s1_write),     //             .write
		.AVS_WriteData   (mm_interconnect_0_piezo_controller_0_s1_writedata), //             .writedata
		.piezo_out       (piezo_controller_piezo_out_export),                 //    piezo_out.export
		.piezo_enable    (piezo_controller_piezo_enable_export),              // piezo_enable.export
		.piezo_enable_in (piezo_controller_piezo_enable_piezo_enable_in),     //             .piezo_enable_in
		.piezo_status    (piezo_controller_piezo_status_export)               // piezo_status.export
	);

	ptp_sync ptp_simple_us_0 (
		.reset                    (rst_controller_reset_out_reset),                             //        reset.reset
		.avalon_slave_address     (mm_interconnect_0_ptp_simple_us_0_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_write       (mm_interconnect_0_ptp_simple_us_0_avalon_slave_write),       //             .write
		.avalon_slave_writedata   (mm_interconnect_0_ptp_simple_us_0_avalon_slave_writedata),   //             .writedata
		.avalon_slave_read        (mm_interconnect_0_ptp_simple_us_0_avalon_slave_read),        //             .read
		.avalon_slave_readdata    (mm_interconnect_0_ptp_simple_us_0_avalon_slave_readdata),    //             .readdata
		.avalon_slave_waitrequest (mm_interconnect_0_ptp_simple_us_0_avalon_slave_waitrequest), //             .waitrequest
		.piezo_interface_in       (ptp_piezo_interface0_piezo_interface_in),                    //  conduit_end.piezo_interface_in
		.piezo_interface_out      (ptp_piezo_interface0_piezo_interface_out),                   //             .piezo_interface_out
		.clock                    (clk_clk)                                                     //        clock.clk
	);

	rtc #(
		.CLOCK_SPEED_HZ (50000000),
		.RTC_RESOLUTION (100)
	) realtime_clock_controll_0 (
		.clock                    (clk_clk),                                                              //   clock_sink.clk
		.event_trigger            (rtc_0_conduit_end_event_trigger),                                      //  conduit_end.event_trigger
		.piezo_enable             (rtc_0_conduit_end_piezo_enable),                                       //             .piezo_enable
		.event_trigger2           (rtc_0_conduit_end_event_trigger2),                                     //             .event_trigger2
		.reset                    (rst_controller_reset_out_reset),                                       //        reset.reset
		.avalon_slave_address     (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_address),     // avalon_slave.address
		.avalon_slave_read        (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_read),        //             .read
		.avalon_slave_readdata    (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_readdata),    //             .readdata
		.avalon_slave_waitrequest (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_waitrequest), //             .waitrequest
		.avalon_slave_write       (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_write),       //             .write
		.avalon_slave_writedata   (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_writedata)    //             .writedata
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                         //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                       //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                        //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                       //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                      //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                       //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                      //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                       //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                      //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                      //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                          //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                        //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                        //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                        //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                       //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                       //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                          //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                        //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                       //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                       //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                         //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                       //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                        //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                       //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                      //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                       //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                      //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                       //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                      //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                      //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                          //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                        //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                        //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                        //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                       //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                       //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                              //                                                     clk_0_clk.clk
		.fpga_key_reset_reset_bridge_in_reset_reset                          (rst_controller_001_reset_out_reset),                                   //                          fpga_key_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                   // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.realtime_clock_controll_0_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                       //         realtime_clock_controll_0_reset_reset_bridge_in_reset.reset
		.fpga_key_s1_address                                                 (mm_interconnect_0_fpga_key_s1_address),                                //                                                   fpga_key_s1.address
		.fpga_key_s1_write                                                   (mm_interconnect_0_fpga_key_s1_write),                                  //                                                              .write
		.fpga_key_s1_readdata                                                (mm_interconnect_0_fpga_key_s1_readdata),                               //                                                              .readdata
		.fpga_key_s1_writedata                                               (mm_interconnect_0_fpga_key_s1_writedata),                              //                                                              .writedata
		.fpga_key_s1_chipselect                                              (mm_interconnect_0_fpga_key_s1_chipselect),                             //                                                              .chipselect
		.fpga_led_s1_address                                                 (mm_interconnect_0_fpga_led_s1_address),                                //                                                   fpga_led_s1.address
		.fpga_led_s1_write                                                   (mm_interconnect_0_fpga_led_s1_write),                                  //                                                              .write
		.fpga_led_s1_readdata                                                (mm_interconnect_0_fpga_led_s1_readdata),                               //                                                              .readdata
		.fpga_led_s1_writedata                                               (mm_interconnect_0_fpga_led_s1_writedata),                              //                                                              .writedata
		.fpga_led_s1_chipselect                                              (mm_interconnect_0_fpga_led_s1_chipselect),                             //                                                              .chipselect
		.id_switch_0_avalon_slave_address                                    (mm_interconnect_0_id_switch_0_avalon_slave_address),                   //                                      id_switch_0_avalon_slave.address
		.id_switch_0_avalon_slave_write                                      (mm_interconnect_0_id_switch_0_avalon_slave_write),                     //                                                              .write
		.id_switch_0_avalon_slave_read                                       (mm_interconnect_0_id_switch_0_avalon_slave_read),                      //                                                              .read
		.id_switch_0_avalon_slave_readdata                                   (mm_interconnect_0_id_switch_0_avalon_slave_readdata),                  //                                                              .readdata
		.id_switch_0_avalon_slave_writedata                                  (mm_interconnect_0_id_switch_0_avalon_slave_writedata),                 //                                                              .writedata
		.id_switch_0_avalon_slave_waitrequest                                (mm_interconnect_0_id_switch_0_avalon_slave_waitrequest),               //                                                              .waitrequest
		.piezo_controller_0_s1_address                                       (mm_interconnect_0_piezo_controller_0_s1_address),                      //                                         piezo_controller_0_s1.address
		.piezo_controller_0_s1_write                                         (mm_interconnect_0_piezo_controller_0_s1_write),                        //                                                              .write
		.piezo_controller_0_s1_read                                          (mm_interconnect_0_piezo_controller_0_s1_read),                         //                                                              .read
		.piezo_controller_0_s1_readdata                                      (mm_interconnect_0_piezo_controller_0_s1_readdata),                     //                                                              .readdata
		.piezo_controller_0_s1_writedata                                     (mm_interconnect_0_piezo_controller_0_s1_writedata),                    //                                                              .writedata
		.ptp_simple_us_0_avalon_slave_address                                (mm_interconnect_0_ptp_simple_us_0_avalon_slave_address),               //                                  ptp_simple_us_0_avalon_slave.address
		.ptp_simple_us_0_avalon_slave_write                                  (mm_interconnect_0_ptp_simple_us_0_avalon_slave_write),                 //                                                              .write
		.ptp_simple_us_0_avalon_slave_read                                   (mm_interconnect_0_ptp_simple_us_0_avalon_slave_read),                  //                                                              .read
		.ptp_simple_us_0_avalon_slave_readdata                               (mm_interconnect_0_ptp_simple_us_0_avalon_slave_readdata),              //                                                              .readdata
		.ptp_simple_us_0_avalon_slave_writedata                              (mm_interconnect_0_ptp_simple_us_0_avalon_slave_writedata),             //                                                              .writedata
		.ptp_simple_us_0_avalon_slave_waitrequest                            (mm_interconnect_0_ptp_simple_us_0_avalon_slave_waitrequest),           //                                                              .waitrequest
		.realtime_clock_controll_0_avalon_slave_address                      (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_address),     //                        realtime_clock_controll_0_avalon_slave.address
		.realtime_clock_controll_0_avalon_slave_write                        (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_write),       //                                                              .write
		.realtime_clock_controll_0_avalon_slave_read                         (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_read),        //                                                              .read
		.realtime_clock_controll_0_avalon_slave_readdata                     (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_readdata),    //                                                              .readdata
		.realtime_clock_controll_0_avalon_slave_writedata                    (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_writedata),   //                                                              .writedata
		.realtime_clock_controll_0_avalon_slave_waitrequest                  (mm_interconnect_0_realtime_clock_controll_0_avalon_slave_waitrequest)  //                                                              .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),             // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
